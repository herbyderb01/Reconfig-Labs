-- read in velocitites, update new position for ball