PLL_25M_inst : PLL_25M PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
